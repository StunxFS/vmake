module vmake

fn test_v_require() {
	require_v('latest')
	require_v('1.2.3')
}

