module main

fn main() {
	// TODO
}

