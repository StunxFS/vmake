module main

// import vmake

fn main() {
	// TODO
}

